//design code given in the question

module top
  (
    input  [1:0]  a,
    output [1:0]  b  
  );
  
assign b = a;
  
  
endmodule
