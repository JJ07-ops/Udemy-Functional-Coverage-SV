//design code given in the question

module top(
  input [1:0] a,b,c,
  output reg [3:0] y
 
);
 
 /*
 User Logic here
 Do not add anything
 ...................
 ..................
 ..................
 ...............
 */
  
endmodule
